LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
	PACKAGE tensorflow_package is
		type padroes is array(0 to 1024) of integer;
		constant bias_mem : padroes := ( -1, others=>0 );
		constant feature_mem : padroes := ( 9, 9, 10, 10, 10, 9, 10, 9, 9, 9, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 7, 7, 9, 9, 9, 10, 10, 10, 10, 10, 10, 9, 9, 9, 10, 10, 10, 10, 10, 10, 9, 9, 9, 8, 8, 8, 9, 9, 9, 8, 8, 8, 7, 7, 9, 9, 9, 10, 10, 10, 10, 10, 10, 10, 9, 9, 10, 10, 10, 10, 10, 9, 9, 7, 6, 6, 6, 7, 7, 8, 8, 8, 8, 8, 8, 7, 9, 9, 10, 10, 10, 10, 10, 10, 10, 10, 10, 11, 11, 9, 10, 10, 9, 9, 6, 6, 6, 5, 5, 4, 5, 5, 7, 8, 8, 8, 8, 7, 9, 9, 10, 10, 10, 10, 10, 10, 10, 10, 10, 15, 12, 9, 9, 8, 6, 4, 5, 7, 7, 6, 6, 5, 4, 5, 5, 6, 8, 8, 8, 8, 9, 8, 8, 9, 10, 10, 10, 10, 10, 10, 10, 11, 9, 8, 6, 4, 4, 4, 5, 7, 7, 7, 7, 5, 6, 5, 3, 4, 6, 8, 8, 8, 7, 6, 2, 5, 9, 10, 10, 10, 10, 10, 10, 9, 8, 7, 6, 4, 4, 4, 5, 8, 9, 7, 6, 6, 7, 5, 3, 2, 4, 8, 8, 8, 8, 6, 2, 4, 8, 10, 10, 10, 10, 10, 8, 7, 8, 9, 7, 5, 5, 5, 4, 7, 10, 8, 6, 6, 6, 5, 3, 3, 3, 6, 8, 8, 10, 6, 3, 7, 9, 10, 10, 10, 10, 10, 7, 7, 9, 9, 7, 5, 5, 5, 5, 5, 8, 9, 7, 5, 5, 5, 4, 3, 2, 4, 8, 8, 11, 8, 5, 9, 10, 9, 9, 9, 12, 14, 12, 9, 10, 9, 7, 5, 5, 4, 3, 4, 8, 8, 8, 6, 5, 5, 5, 4, 3, 2, 5, 8, 11, 6, 8, 10, 11, 9, 9, 7, 13, 14, 13, 10, 11, 9, 7, 7, 4, 5, 2, 5, 10, 9, 9, 6, 5, 6, 5, 4, 3, 2, 3, 6, 11, 6, 8, 10, 11, 10, 10, 8, 7, 12, 12, 10, 11, 11, 8, 7, 6, 5, 2, 7, 13, 10, 9, 5, 5, 5, 6, 5, 4, 3, 3, 4, 11, 5, 7, 10, 10, 10, 11, 9, 6, 10, 10, 8, 11, 13, 10, 7, 7, 7, 3, 9, 12, 9, 7, 5, 5, 5, 5, 5, 5, 4, 4, 4, 11, 5, 9, 11, 7, 8, 10, 10, 6, 9, 9, 10, 11, 14, 11, 8, 7, 7, 4, 9, 11, 9, 7, 5, 5, 4, 5, 6, 6, 5, 6, 5, 12, 6, 10, 11, 6, 6, 9, 10, 6, 7, 8, 12, 11, 10, 9, 9, 9, 6, 4, 9, 11, 8, 8, 6, 5, 5, 5, 6, 7, 6, 6, 7, 12, 8, 10, 11, 8, 4, 8, 9, 7, 8, 8, 14, 15, 9, 8, 8, 7, 6, 5, 9, 10, 9, 7, 5, 4, 5, 6, 7, 7, 6, 7, 8, 12, 9, 10, 11, 10, 4, 7, 8, 8, 6, 9, 10, 10, 8, 7, 7, 6, 6, 7, 10, 9, 9, 8, 6, 4, 4, 5, 6, 6, 7, 9, 9, 13, 10, 10, 11, 11, 5, 6, 9, 9, 6, 8, 7, 7, 7, 6, 7, 5, 6, 9, 7, 4, 8, 8, 4, 3, 3, 4, 6, 7, 8, 9, 8, 13, 11, 10, 10, 11, 7, 5, 8, 9, 8, 6, 4, 8, 7, 8, 9, 5, 5, 9, 8, 7, 6, 4, 4, 2, 4, 5, 8, 9, 10, 9, 9, 12, 11, 10, 10, 11, 9, 5, 7, 7, 8, 9, 4, 8, 6, 9, 11, 7, 4, 8, 8, 8, 5, 3, 3, 2, 5, 7, 10, 10, 10, 9, 9, 10, 12, 11, 11, 11, 9, 6, 8, 10, 6, 5, 5, 5, 7, 11, 11, 9, 6, 5, 5, 3, 2, 2, 1, 2, 3, 6, 9, 9, 8, 7, 7, 7, 12, 11, 11, 11, 8, 5, 9, 15, 13, 8, 8, 9, 11, 11, 12, 10, 7, 6, 3, 2, 2, 3, 3, 3, 3, 4, 4, 4, 4, 3, 3, 4, 10, 10, 11, 11, 8, 6, 13, 15, 15, 13, 7, 7, 7, 7, 7, 6, 4, 4, 3, 3, 3, 3, 3, 3, 3, 2, 3, 3, 3, 2, 2, 2, 6, 9, 10, 11, 10, 10, 15, 15, 14, 6, 3, 3, 3, 3, 3, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 3, 3, 3, 3, 2, 1, 1, 3, 8, 10, 8, 12, 15, 15, 8, 3, 3, 3, 3, 3, 3, 2, 2, 2, 2, 2, 2, 2, 2, 2, 3, 3, 3, 3, 3, 2, 3, 3, 1, 2, 4, 8, 8, 13, 16, 11, 4, 3, 3, 3, 3, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 3, 3, 4, 3, 3, 3, 4, 5, 3, 2, 1, 2, 4, 8, 14, 15, 7, 3, 3, 3, 3, 2, 2, 2, 2, 2, 2, 2, 2, 2, 3, 3, 3, 2, 2, 2, 3, 4, 5, 4, 3, 2, 1, 2, 2, 4, 12, 13, 6, 4, 3, 3, 3, 3, 2, 2, 2, 3, 2, 2, 3, 2, 2, 3, 2, 2, 1, 2, 4, 4, 2, 3, 3, 2, 2, 2, 2, 2, 6, 10, 4, 3, 3, 3, 3, 3, 3, 2, 2, 2, 2, 3, 2, 2, 2, 2, 2, 2, 2, 3, 2, 1, 0, 3, 4, 2, 1, 2, 2, 2, 2, 4, 3, 1, 1, 2, 3, 3, 3, 3, 3, 3, 3, 3, 3, 2, 2, 2, 2, 3, 4, 4, 3, 2, 0, 2, 3, 3, 2, 2, 2, 2, 2, 2, 2, 1, 1, 1, 1, 1, 2, 2, 3, 3, 4, 4, 4, 3, 2, 2, 3, 5, 6, 5, 3, 1, 1, 1, 3, 3, 2, 2, 2, 2, 2, 2, 2, 1, 1, 1, 1, 1, 1, 1, 2, 2, 3, 4, 4, 3, 3, 2, 4, 5, 6, 5, 3, 1, 2, 1, others=>0 );
		constant weight_mem : padroes := ( 4, 1, -2, 2, 0, -5, -2, 0, -5, others=>0 );
		constant gold : padroes := ( 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, others=>0 );
END tensorflow_package;
